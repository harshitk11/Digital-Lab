`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:42:18 09/30/2016 
// Design Name: 
// Module Name:    index_mem 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module index_mem(i1,i2,cnt1,cnt2,r1,r2);
input i1,i2,cnt1,cnt2;
output r1,r2;
wire [3:0]	i1,i2,cnt1,cnt2;
reg [3:0] r1,r2;




endmodule
